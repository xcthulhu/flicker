../lfsr_tb.vhdl